�� sr java.util.ArrayListx����a� I sizexp   w   sr +jlhthdfinalboardgame.boardmanagement.Player񷶩���� I scoreL colort )Ljlhthdfinalboardgame/table/PlayerColors;L remainingBeadst Ljava/lang/Integer;[ 
scoreArrayt ([Ljlhthdfinalboardgame/table/BeadColors;L selectedColort 'Ljlhthdfinalboardgame/table/BeadColors;L startingBeadsq ~ xp    ~r 'jlhthdfinalboardgame.table.PlayerColors          xr java.lang.Enum          xpt WHITEsr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   ur ([Ljlhthdfinalboardgame.table.BeadColors;�.3�L�M�  xp   ~r %jlhthdfinalboardgame.table.BeadColors          xq ~ 	t BLUE~q ~ t GREEN~q ~ t RED~q ~ t YELLOWq ~ sq ~    sq ~     ~q ~ t BLACKsq ~    uq ~    q ~ q ~ q ~ q ~ q ~ q ~ xq ~ ~r 7jlhthdfinalboardgame.boardmanagement.BoardManager$Phase          xq ~ 	t COLORw   sr  jlhthdfinalboardgame.table.Table�d&�E I numColsI numRowsL tablet Ljava/util/ArrayList;xp      sq ~     w   sq ~     w   sr ,jlhthdfinalboardgame.table.PlayerColorObject(Lz4w� L colorq ~ xp~q ~ t NONEsq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ 
sq ~ (q ~ sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ 
sq ~ (q ~ 
sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *xsq ~     w   sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *sq ~ (q ~ *xxsq ~ #      	sq ~     	w   	sq ~     w   sr *jlhthdfinalboardgame.table.BeadColorObject�2Bct�� L colorq ~ xp~q ~ t NONEsq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ sq ~ ]q ~ sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xsq ~     w   sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _sq ~ ]q ~ _xx